module	testbench();
reg clk,rst,rx;
wire tx;
top test(.clk(clk),.rst(rst),.rx(rx),.tx(tx));
initial
begin
    rst = 1;
    #50000 rst = 0;
    #20000000 $stop;
end
initial
begin
    clk = 0;
    forever #1 clk = ~clk;
end
initial
begin
    //在rst重置后，再加上一堆空闲帧 
    //每一帧以866开始（0），8个1736数据位，再以866（0）结束
    rx = 0;
    #100000      rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 0

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 2

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 3

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 4

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 5

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 6

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 7

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 8

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 9

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 10

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 11

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 12

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 13

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 14

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 15

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 16

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 17

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 18

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 19

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 20

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 21

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 22

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 23

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 24

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 25

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 26

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 27

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 28

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 29

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 30

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 31

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 32

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 33

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 34

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 35

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 36

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 37

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 38

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 39

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 40

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 41

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 42

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 43

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 44

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 45

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 46

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 47

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 48

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 49

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 50

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 51

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 52

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 53

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 54

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 55

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 56

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 57

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 58

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 59

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 60

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 61

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 62

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 63

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 64

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 65

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 66

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 67

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 68

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 69

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 70

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 71

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 72

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 73

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 74

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 75

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 76

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 77

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 78

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 79

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 80

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 81

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 82

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 83

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 84

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 85

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 86

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 87

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 88

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 89

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 90

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 91

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 92

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 93

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 94

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 95

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 96

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 97

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 98

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 99

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 100

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 101

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 102

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 103

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 104

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 105

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 106

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 107

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 108

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 109

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 110

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 111

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 112

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 113

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 114

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 115

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 116

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 117

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 118

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 119

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 120

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 121

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 122

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 123

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 124

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 125

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 126

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 127

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 128

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 129

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 130

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 131

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 132

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 133

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 134

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 135

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 136

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 137

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 138

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 139

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 140

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 141

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 142

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 143

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 144

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 145

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 146

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 147

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 148

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 149

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 150

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 151

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 152

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 153

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 154

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 155

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 156

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 157

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 158

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 159

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 160

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 161

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 162

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 163

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 164

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 165

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 166

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 167

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 168

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 169

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 170

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 171

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 172

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 173

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 174

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 175

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 176

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 177

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 178

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 179

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 180

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 181

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 182

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 183

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 184

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 185

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 186

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 187

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 188

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 189

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 190

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 191

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 192

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 193

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 194

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 195

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 196

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 197

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 198

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 199

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 200

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 201

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 202

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 203

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 204

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 205

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 206

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 207

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 208

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 209

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 210

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 211

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 212

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 213

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 214

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 215

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 216

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 217

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 218

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 219

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 220

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 221

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 222

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 223

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 224

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 225

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 226

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 227

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 228

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 229

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 230

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 231

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 232

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 233

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 234

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 235

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 236

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 237

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 238

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 239

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 240

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 241

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 242

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 243

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 244

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 245

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 246

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 247

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 248

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 249

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 250

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 251

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 252

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 253

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 254

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 255

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 256

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 257

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 258

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 259

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 260

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 261

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 262

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 263

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 264

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 265

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 266

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 267

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 268

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 269

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 270

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 271

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 272

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 273

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 274

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 275

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 276

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 277

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 278

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 279

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 280

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 281

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 282

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 283

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 284

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 285

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 286

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 287

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 288

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 289

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 290

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 291

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 292

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 293

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 294

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 295

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 296

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 297

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 298

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 299

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 300

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 301

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 302

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 303

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 304

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 305

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 306

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 307

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 308

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 309

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 310

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 311

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 312

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 313

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 314

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 315

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 316

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 317

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 318

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 319

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 320

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 321

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 322

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 323

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 324

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 325

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 326

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 327

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 328

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 329

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 330

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 331

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 332

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 333

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 334

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 335

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 336

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 337

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 338

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 339

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 340

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 341

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 342

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 343

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 344

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 345

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 346

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 347

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 348

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 349

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 350

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 351

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 352

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 353

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 354

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 355

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 356

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 357

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 358

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 359

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 360

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 361

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 362

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 363

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 364

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 365

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 366

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 367

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 368

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 369

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 370

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 371

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 372

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 373

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 374

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 375

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 376

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 377

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 378

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 379

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 380

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 381

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 382

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 383

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 384

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 385

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 386

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 387

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 388

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 389

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 390

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 391

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 392

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 393

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 394

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 395

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 396

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 397

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 398

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 399

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 400

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 401

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 402

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 403

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 404

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 405

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 406

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 407

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 408

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 409

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 410

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 411

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 412

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 413

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 414

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 415

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 416

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 417

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 418

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 419

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 420

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 421

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 422

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 423

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 424

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 425

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 426

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 427

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 428

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 429

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 430

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 431

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 432

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 433

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 434

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 435

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 436

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 437

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 438

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 439

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 440

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 441

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 442

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 443

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 444

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 445

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 446

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 447

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 448

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 449

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 450

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 451

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 452

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 453

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 454

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 455

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 456

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 457

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 458

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 459

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 460

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 461

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 462

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 463

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 464

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 465

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 466

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 467

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 468

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 469

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 470

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 471

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 472

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 473

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 474

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 475

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 476

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 477

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 478

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 479

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 480

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 481

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 482

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 483

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 484

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 485

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 486

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 487

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 488

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 489

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 490

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 491

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 492

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 493

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 494

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 495

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 496

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 497

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 498

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 499

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 500

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 501

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 502

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 503

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 504

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 505

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 506

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 507

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 508

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 509

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 510

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 511

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 512

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 513

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 514

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 515

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 516

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 517

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 518

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 519

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 520

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 521

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 522

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 523

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 524

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 525

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 526

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 527

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 528

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 529

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 530

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 531

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 532

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 533

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 534

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 535

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 536

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 537

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 538

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 539

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 540

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 541

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 542

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 543

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 544

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 545

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 546

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 547

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 548

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 549

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 550

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 551

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 552

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 553

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 554

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 555

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 556

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 557

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 558

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 559

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 560

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 561

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 562

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 563

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 564

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 565

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 566

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 567

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 568

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 569

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 570

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 571

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 572

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 573

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 574

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 575

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 576

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 577

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 578

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 579

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 580

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 581

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 582

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 583

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 584

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 585

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 586

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 587

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 588

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 589

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 590

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 591

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 592

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 593

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 594

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 595

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 596

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 597

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 598

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 599

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 600

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 601

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 602

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 603

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 604

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 605

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 606

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 607

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 608

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 609

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 610

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 611

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 612

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 613

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 614

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 615

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 616

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 617

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 618

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 619

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 620

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 621

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 622

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 623

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 624

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 625

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 626

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 627

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 628

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 629

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 630

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 631

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 632

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 633

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 634

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 635

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 636

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 637

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 638

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 639

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 640

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 641

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 642

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 643

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 644

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 645

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 646

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 647

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 648

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 649

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 650

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 651

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 652

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 653

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 654

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 655

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 656

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 657

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 658

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 659

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 660

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 661

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 662

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 663

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 664

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 665

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 666

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 667

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 668

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 669

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 670

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 671

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 672

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 673

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 674

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 675

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 676

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 677

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 678

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 679

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 680

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 681

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 682

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 683

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 684

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 685

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 686

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 687

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 688

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 689

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 690

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 691

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 692

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 693

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 694

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 695

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 696

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 697

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 698

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 699

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 700

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 701

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 702

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 703

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 704

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 705

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 706

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 707

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 708

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 709

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 710

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 711

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 712

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 713

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 714

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 715

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 716

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 717

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 718

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 719

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 720

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 721

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 722

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 723

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 724

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 725

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 726

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 727

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 728

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 729

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 730

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 731

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 732

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 733

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 734

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 735

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 736

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 737

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 738

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 739

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 740

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 741

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 742

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 743

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 744

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 745

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 746

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 747

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 748

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 749

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 750

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 751

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 752

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 753

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 754

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 755

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 756

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 757

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 758

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 759

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 760

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 761

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 762

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 763

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 764

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 765

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 766

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 767

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 768

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 769

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 770

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 771

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 772

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 773

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 774

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 775

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 776

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 777

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 778

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 779

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 780

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 781

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 782

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 783

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 784

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 785

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 786

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 787

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 788

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 789

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 790

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 791

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 792

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 793

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 794

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 795

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 796

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 797

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 798

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 799

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 800

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 801

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 802

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 803

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 804

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 805

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 806

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 807

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 808

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 809

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 810

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 811

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 812

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 813

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 814

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 815

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 816

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 817

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 818

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 819

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 820

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 821

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 822

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 823

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 824

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 825

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 826

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 827

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 828

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 829

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 830

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 831

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 832

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 833

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 834

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 835

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 836

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 837

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 838

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 839

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 840

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 841

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 842

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 843

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 844

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 845

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 846

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 847

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 848

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 849

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 850

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 851

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 852

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 853

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 854

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 855

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 856

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 857

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 858

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 859

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 860

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 861

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 862

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 863

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 864

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 865

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 866

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 867

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 868

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 869

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 870

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 871

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 872

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 873

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 874

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 875

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 876

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 877

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 878

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 879

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 880

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 881

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 882

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 883

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 884

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 885

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 886

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 887

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 888

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 889

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 890

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 891

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 892

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 893

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 894

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 895

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 896

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 897

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 898

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 899

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 900

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 901

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 902

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 903

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 904

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 905

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 906

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 907

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 908

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 909

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 910

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 911

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 912

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 913

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 914

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 915

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 916

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 917

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 918

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 919

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 920

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 921

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #866        rx = 0;
//num == 922

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 923

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 924

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 925

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 926

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 927

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 928

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 929

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 930

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 931

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 932

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 933

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 934

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 935

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 936

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 937

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 938

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 939

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 940

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 941

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 942

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 943

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 944

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 945

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 946

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 947

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 948

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 949

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 950

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 951

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 952

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 953

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 954

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 955

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 956

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 957

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 958

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 959

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 960

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 961

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 962

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 963

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 964

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 965

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 966

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 967

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 968

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 969

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 970

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 971

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 972

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 973

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 974

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 975

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 976

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 977

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 978

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 979

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 980

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 981

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 982

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 983

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 984

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 985

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 986

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 987

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 988

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 989

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 990

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 991

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 992

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 993

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 994

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 995

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 996

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 997

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 998

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 999

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1000

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1001

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1002

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1003

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1004

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1005

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1006

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1007

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1008

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1009

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1010

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1011

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1012

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1013

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1014

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1015

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1016

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1017

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1018

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1019

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1020

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1021

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1022

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1023

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1024

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1025

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1026

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1027

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1028

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1029

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1030

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1031

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1032

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1033

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1034

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1035

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1036

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1037

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1038

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1039

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1040

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1041

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1042

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1043

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1044

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1045

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1046

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1047

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1048

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1049

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1050

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1051

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1052

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1053

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1054

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1055

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1056

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1057

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1058

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1059

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1060

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1061

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1062

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1063

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1064

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1065

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1066

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1067

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1068

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1069

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1070

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1071

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1072

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1073

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1074

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1075

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1076

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1077

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1078

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1079

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1080

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1081

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1082

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1083

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1084

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1085

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1086

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1087

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1088

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1089

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1090

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1091

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1092

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1093

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1094

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1095

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1096

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1097

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1098

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1099

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1100

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1101

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1102

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1103

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1104

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1105

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1106

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1107

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1108

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1109

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1110

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1111

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1112

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1113

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1114

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1115

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1116

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1117

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1118

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1119

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1120

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1121

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1122

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1123

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1124

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1125

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1126

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1127

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1128

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1129

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1130

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1131

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1132

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1133

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1134

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1135

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1136

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1137

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1138

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1139

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1140

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1141

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1142

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1143

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1144

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1145

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1146

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1147

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1148

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1149

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1150

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1151

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1152

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1153

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1154

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1155

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1156

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1157

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1158

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1159

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1160

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1161

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1162

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1163

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1164

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1165

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1166

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1167

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1168

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1169

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1170

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1171

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1172

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1173

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1174

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1175

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1176

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1177

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1178

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1179

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1180

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1181

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1182

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1183

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1184

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1185

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1186

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1187

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1188

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1189

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1190

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1191

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1192

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1193

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1194

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1195

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1196

    #866        rx = 0;
    #866        rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1197

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1198

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
//num == 1199

    #866        rx = 0;
    #866        rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #866        rx = 0;
end
endmodule
