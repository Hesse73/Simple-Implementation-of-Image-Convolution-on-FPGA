module	testbench();
reg clk,rst,rx;
wire tx;
top test(.clk(clk),.rst(rst),.rx(rx),.tx(tx));
initial
begin
    rst = 1;
    #50000 rst = 0;
    #20000000 $stop;
end
initial
begin
    clk = 0;
    forever #1 clk = ~clk;
end
initial
begin
    //每一帧以866开始（0），8个1736数据位，再以866（0）结束
    rx = 0;
    #100000      rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 0

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 2

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 3

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 4

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 5

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 6

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 7

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 8

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 9

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 10

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 11

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 12

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 13

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 14

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 15

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 16

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 17

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 18

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 19

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 20

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 21

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 22

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 23

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 24

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 25

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 26

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 27

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 28

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 29

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 30

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 31

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 32

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 33

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 34

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 35

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 36

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 37

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 38

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 39

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 40

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 41

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 42

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 43

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 44

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 45

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 46

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 47

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 48

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 49

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 50

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 51

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 52

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 53

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 54

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 55

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 56

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 57

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 58

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 59

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 60

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 61

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 62

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 63

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 64

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 65

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 66

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 67

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 68

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 69

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 70

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 71

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 72

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 73

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 74

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 75

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 76

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 77

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 78

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 79

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 80

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 81

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 82

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 83

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 84

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 85

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 86

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 87

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 88

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 89

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 90

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 91

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 92

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 93

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 94

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 95

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 96

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 97

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 98

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 99

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 100

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 101

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 102

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 103

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 104

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 105

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 106

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 107

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 108

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 109

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 110

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 111

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 112

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 113

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 114

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 115

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 116

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 117

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 118

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 119

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 120

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 121

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 122

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 123

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 124

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 125

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 126

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 127

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 128

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 129

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 130

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 131

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 132

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 133

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 134

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 135

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 136

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 137

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 138

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 139

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 140

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 141

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 142

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 143

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 144

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 145

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 146

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 147

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 148

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 149

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 150

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 151

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 152

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 153

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 154

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 155

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 156

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 157

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 158

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 159

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 160

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 161

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 162

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 163

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 164

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 165

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 166

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 167

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 168

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 169

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 170

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 171

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 172

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 173

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 174

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 175

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 176

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 177

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 178

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 179

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 180

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 181

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 182

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 183

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 184

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 185

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 186

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 187

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 188

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 189

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 190

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 191

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 192

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 193

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 194

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 195

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 196

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 197

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 198

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 199

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 200

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 201

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 202

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 203

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 204

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 205

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 206

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 207

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 208

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 209

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 210

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 211

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 212

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 213

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 214

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 215

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 216

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 217

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 218

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 219

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 220

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 221

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 222

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 223

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 224

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 225

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 226

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 227

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 228

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 229

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 230

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 231

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 232

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 233

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 234

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 235

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 236

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 237

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 238

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 239

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 240

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 241

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 242

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 243

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 244

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 245

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 246

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 247

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 248

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 249

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 250

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 251

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 252

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 253

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 254

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 255

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 256

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 257

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 258

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 259

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 260

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 261

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 262

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 263

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 264

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 265

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 266

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 267

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 268

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 269

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 270

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 271

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 272

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 273

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 274

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 275

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 276

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 277

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 278

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 279

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 280

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 281

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 282

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 283

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 284

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 285

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 286

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 287

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 288

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 289

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 290

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 291

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 292

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 293

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 294

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 295

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 296

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 297

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 298

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 299

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 300

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 301

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 302

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 303

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 304

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 305

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 306

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 307

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 308

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 309

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 310

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 311

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 312

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 313

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 314

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 315

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 316

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 317

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 318

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 319

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 320

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 321

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 322

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 323

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 324

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 325

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 326

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 327

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 328

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 329

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 330

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 331

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 332

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 333

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 334

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 335

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 336

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 337

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 338

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 339

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 340

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 341

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 342

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 343

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 344

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 345

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 346

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 347

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 348

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 349

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 350

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 351

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 352

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 353

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 354

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 355

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 356

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 357

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 358

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 359

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 360

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 361

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 362

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 363

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 364

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 365

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 366

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 367

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 368

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 369

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 370

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 371

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 372

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 373

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 374

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 375

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 376

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 377

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 378

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 379

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 380

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 381

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 382

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 383

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 384

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 385

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 386

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 387

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 388

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 389

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 390

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 391

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 392

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 393

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 394

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 395

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 396

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 397

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 398

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 399

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 400

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 401

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 402

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 403

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 404

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 405

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 406

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 407

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 408

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 409

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 410

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 411

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 412

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 413

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 414

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 415

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 416

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 417

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 418

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 419

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 420

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 421

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 422

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 423

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 424

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 425

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 426

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 427

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 428

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 429

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 430

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 431

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 432

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 433

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 434

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 435

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 436

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 437

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 438

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 439

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 440

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 441

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 442

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 443

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 444

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 445

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 446

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 447

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 448

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 449

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 450

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 451

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 452

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 453

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 454

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 455

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 456

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 457

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 458

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 459

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 460

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 461

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 462

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 463

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 464

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 465

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 466

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 467

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 468

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 469

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 470

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 471

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 472

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 473

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 474

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 475

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 476

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 477

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 478

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 479

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 480

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 481

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 482

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 483

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 484

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 485

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 486

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 487

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 488

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 489

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 490

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 491

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 492

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 493

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 494

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 495

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 496

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 497

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 498

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 499

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 500

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 501

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 502

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 503

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 504

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 505

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 506

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 507

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 508

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 509

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 510

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 511

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 512

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 513

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 514

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 515

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 516

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 517

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 518

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 519

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 520

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 521

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 522

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 523

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 524

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 525

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 526

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 527

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 528

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 529

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 530

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 531

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 532

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 533

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 534

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 535

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 536

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 537

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 538

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 539

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 540

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 541

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 542

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 543

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 544

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 545

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 546

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 547

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 548

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 549

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 550

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 551

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 552

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 553

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 554

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 555

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 556

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 557

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 558

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 559

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 560

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 561

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 562

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 563

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 564

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 565

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 566

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 567

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 568

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 569

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 570

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 571

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 572

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 573

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 574

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 575

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 576

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 577

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 578

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 579

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 580

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 581

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 582

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 583

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 584

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 585

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 586

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 587

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 588

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 589

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 590

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 591

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 592

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 593

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 594

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 595

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 596

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 597

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 598

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 599

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 600

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 601

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 602

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 603

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 604

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 605

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 606

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 607

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 608

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 609

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 610

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 611

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 612

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 613

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 614

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 615

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 616

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 617

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 618

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 619

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 620

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 621

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 622

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 623

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 624

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 625

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 626

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 627

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 628

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 629

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 630

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 631

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 632

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 633

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 634

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 635

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 636

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 637

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 638

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 639

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 640

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 641

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 642

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 643

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 644

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 645

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 646

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 647

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 648

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 649

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 650

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 651

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 652

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 653

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 654

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 655

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 656

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 657

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 658

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 659

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 660

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 661

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 662

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 663

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 664

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 665

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 666

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 667

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 668

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 669

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 670

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 671

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 672

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 673

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 674

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 675

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 676

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 677

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 678

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 679

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 680

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 681

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 682

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 683

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 684

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 685

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 686

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 687

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 688

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 689

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 690

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 691

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 692

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 693

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 694

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 695

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 696

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 697

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 698

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 699

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 700

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 701

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 702

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 703

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 704

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 705

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 706

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 707

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 708

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 709

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 710

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 711

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 712

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 713

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 714

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 715

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 716

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 717

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 718

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 719

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 720

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 721

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 722

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 723

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 724

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 725

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 726

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 727

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 728

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 729

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 730

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 731

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 732

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 733

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 734

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 735

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 736

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 737

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 738

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 739

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 740

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 741

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 742

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 743

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 744

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 745

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 746

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 747

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 748

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 749

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 750

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 751

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 752

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 753

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 754

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 755

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 756

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 757

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 758

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 759

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 760

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 761

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 762

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 763

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 764

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 765

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 766

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 767

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 768

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 769

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 770

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 771

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 772

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 773

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 774

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 775

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 776

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 777

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 778

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 779

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 780

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 781

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 782

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 783

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 784

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 785

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 786

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 787

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 788

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 789

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 790

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 791

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 792

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 793

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 794

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 795

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 796

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 797

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 798

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 799

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 800

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 801

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 802

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 803

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 804

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 805

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 806

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 807

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 808

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 809

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 810

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 811

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 812

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 813

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 814

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 815

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 816

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 817

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 818

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 819

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 820

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 821

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 822

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 823

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 824

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 825

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 826

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 827

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 828

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 829

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 830

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 831

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 832

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 833

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 834

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 835

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 836

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 837

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 838

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 839

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 840

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 841

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 842

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 843

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 844

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 845

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 846

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 847

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 848

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 849

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 850

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 851

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 852

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 853

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 854

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 855

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 856

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 857

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 858

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 859

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 860

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 861

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 862

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 863

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 864

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 865

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 866

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 867

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 868

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 869

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 870

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 871

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 872

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 873

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 874

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 875

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 876

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 877

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 878

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 879

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 880

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 881

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 882

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 883

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 884

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 885

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 886

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 887

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 888

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 889

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 890

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 891

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 892

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 893

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 894

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 895

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 896

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 897

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 898

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 899

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 900

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 901

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 902

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 903

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 904

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 905

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 906

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 907

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 908

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 909

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 910

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 911

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 912

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 913

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 914

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 915

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 916

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 917

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 918

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 919

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 920

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 921

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 922

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 923

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 924

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 925

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 926

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 927

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 928

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 929

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 930

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 931

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 932

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 933

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 934

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 935

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 936

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 937

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 938

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 939

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 940

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 941

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 942

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 943

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 944

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 945

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 946

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 947

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 948

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 949

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 950

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 951

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 952

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 953

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 954

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 955

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 956

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 957

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 958

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 959

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 960

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 961

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 962

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 963

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 964

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 965

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 966

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 967

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 968

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 969

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 970

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 971

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 972

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 973

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 974

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 975

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 976

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 977

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 978

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 979

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 980

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 981

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 982

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 983

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 984

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 985

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 986

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 987

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 988

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 989

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 990

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 991

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 992

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 993

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 994

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 995

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 996

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 997

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 998

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 999

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1000

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1001

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1002

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1003

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1004

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1005

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1006

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1007

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1008

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1009

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1010

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1011

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1012

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1013

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1014

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1015

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1016

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1017

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1018

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1019

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1020

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1021

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1022

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1023

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1024

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1025

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1026

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1027

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1028

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1029

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1030

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1031

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1032

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1033

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1034

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1035

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1036

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1037

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1038

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1039

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1040

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1041

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1042

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1043

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1044

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1045

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1046

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1047

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1048

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1049

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1050

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1051

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1052

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1053

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1054

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1055

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1056

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1057

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1058

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1059

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1060

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1061

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1062

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1063

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1064

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1065

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1066

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1067

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1068

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1069

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1070

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1071

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1072

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1073

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1074

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1075

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1076

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1077

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1078

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1079

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1080

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1081

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1082

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1083

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1084

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1085

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1086

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1087

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1088

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1089

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1090

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1091

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1092

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1093

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1094

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1095

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1096

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1097

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1098

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1099

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1100

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1101

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1102

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1103

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1104

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1105

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1106

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1107

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1108

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1109

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1110

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1111

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1112

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1113

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1114

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1115

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1116

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1117

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1118

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1119

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1120

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1121

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1122

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1123

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1124

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1125

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1126

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1127

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1128

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1129

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1130

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1131

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1132

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1133

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1134

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1135

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1136

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1137

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1138

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1139

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1140

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1141

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1142

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1143

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1144

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1145

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1146

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1147

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1148

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1149

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1150

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1151

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1152

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1153

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1154

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1155

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1156

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1157

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1158

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1159

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1160

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1161

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1162

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1163

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1164

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1165

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1166

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1167

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1168

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1169

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1170

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1171

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1172

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1173

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1174

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1175

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1176

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1177

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1178

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1179

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1180

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1181

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1182

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1183

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1184

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1185

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1186

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1187

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1188

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1189

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1190

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1191

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1192

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1193

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1194

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1195

    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1196

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1197

    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1198

    #1736       rx = 1;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
 //num = 1199

    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 0;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 1;
    #1736       rx = 0;
    #1736        rx = 0;
end
endmodule
